/**********************************************************
 Start Date: 11 Sept 2015
 Finish Date: 11 Sept 2015
 Author: Mayur Kubavat
 
 Module: Test Package
 Filename: test_pkg.sv
**********************************************************/

package ahb_test_pkg;

        `include "uvm_macros.svh"
        import uvm_pkg::*;

        `include "tb_defs.svh"


        `include "ahb_mxtn.svh"
        `include "ahb_sxtn.svh"

        `include "ahb_magent_config.svh"
        `include "ahb_mseqr.svh"
        `include "ahb_mdriver.svh"
        `include "ahb_mmonitor.svh"

        `include "ahb_sagent_config.svh"
        `include "ahb_sseqr.svh"
        `include "ahb_sdriver.svh"
        `include "ahb_smonitor.svh"

        `include "reset_seqr.svh"
        `include "reset_driver.svh"

        `include "env_config.svh"
        `include "ahb_vseqr.svh"
        `include "reset_agent.svh"
        `include "ahb_magent.svh"
        `include "ahb_sagent.svh"
        `include "ahb_coverage.svh"

        `include "ahb_env.svh"

        `include "reset_seqs.svh"
        `include "ahb_mseqs.svh"
        `include "ahb_sseqs.svh"
        `include "ahb_vseqs.svh"

        `include "ahb_test.svh"

endpackage

